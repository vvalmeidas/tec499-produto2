//------------------------------------------------------------------------------
//	Module:	FPGA_TOP_MIV
//	Desc:	Top level interface from a Mercurio FPGA board
//------------------------------------------------------------------------------

module LCD_Controller_TOP
	(
		//------------------------------------------------------------------
		//	Clock & Reset Inputs
		//------------------------------------------------------------------
		Clock,
		Reset,
		//------------------------------------------------------------------
		
		//------------------------------------------------------------------
		//	Inputs
		//------------------------------------------------------------------
		//------------------------------------------------------------------
		
		//------------------------------------------------------------------
		//	Outputs
		//------------------------------------------------------------------
		Estado,
		Enable,
		RS,
		RW,
		Dados
		//------------------------------------------------------------------
	);

	////////////////////////	Clock Input	 	////////////////////////
	input			Clock;						
	////////////////////////	RGB LED		   ////////////////////////
	output			[2:0] Estado;							//	RGB LED Green

	wire	[2:0]				estado_inicializador;
	wire			 	Enable;
	output				RS;
	output				RW;
	output	[7:0]		Dados;

	//--------------------------------------------------------------------------
	//	Parameters
	//--------------------------------------------------------------------------
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Parse input from buttons
	//--------------------------------------------------------------------------

	Inicializador_LCD	Instancia_Inicializador	(	
						.Clock(				Clock),
						.Reset(				Reset),
						.Estado(				estado_inicializador),
						.Enable(				Enter)),
						.RS(				Enter)),
						.RW(				Enter)),
						.Dados(				Enter));

						

	Lab2Lock		Lab2LockFSM (
						.Clock(				clock_50MHz),
						.Reset(				LockReset),
						.Enter(				Enter),
						.Digit(				Digit),
						.State(				State),
						.Open(				Open),
						.Fail(				Fail));
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Output Logic
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------	

endmodule